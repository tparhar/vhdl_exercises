library IEEE; use IEEE.STD_LOGIC_1164.all;

entity generic_rca is
	generic(N: integer := 4);
	port(cin:  in STD_LOGIC;
			 a, b: in STD_LOGIC_VECTOR(N-1 downto 0);
			 cout: out STD_LOGIC;
			 s:    out STD_LOGIC_VECTOR(N-1 downto 0));
end generic_rca;

architecture struct of generic_rca is
	component fulladder
		port(a, b, cin: in STD_LOGIC;
				 s, cout: 	out STD_LOGIC);
	end component;
	signal carry_sig: STD_LOGIC_VECTOR(N-1 downto 0);
	signal carry_in:  STD_LOGIC_VECTOR(N-1 downto 0);
begin

	-- initialize carry_in to be cin, and follow carry out by shifting to the left one bit each time
	-- carry out changes
	carry_in <= (carry_sig(N-2 downto 0) & cin);
	
	Adders:
	for i in 0 to N-1 generate
		begin
		ADD1:
				fulladder port map(
						a => a(i),
						b => b(i),
						cin => carry_in(i),
						s => s(i),
						cout => carry_sig(i)
				);
		end generate;
		
		Carry_Out:
				cout <= carry_sig(N-1);
end struct;