library IEEE; use IEEE.STD_LOGIC_1164.all;

entity blockgates is
	port(a, b: 																						 in STD_LOGIC;
			 y_not, y_and, y_or, y_xor, y_nand, y_nor, y_xnor: out STD_LOGIC);
end blockgates;

architecture behv of blockgates is
begin
	y_not <= not a;
	y_and <= a and b;
	y_or <= a or b;
	y_xor <= a xor b;
	y_nand <= a nand b;
	y_nor <= a nor b;
	y_xnor <= a xnor b;
end behv;